package cntr_operations;

  typedef enum { cntr_op_state_1, cntr_op_state_2, cntr_op_state_3 } cntr_operations_t;

endpackage